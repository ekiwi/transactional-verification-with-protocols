module BrCondArea(
  input  [31:0] io_rs1,
  input  [31:0] io_rs2,
  input  [2:0]  io_br_type,
  output        io_taken
);
  wire [31:0] diff; // @[BrCond.scala 37:21]
  wire  neq; // @[BrCond.scala 38:19]
  wire  eq; // @[BrCond.scala 39:14]
  wire  _T_1; // @[BrCond.scala 40:26]
  wire  _T_2; // @[BrCond.scala 40:45]
  wire  isSameSign; // @[BrCond.scala 40:35]
  wire  _T_3; // @[BrCond.scala 41:34]
  wire  lt; // @[BrCond.scala 41:17]
  wire  ltu; // @[BrCond.scala 42:17]
  wire  ge; // @[BrCond.scala 43:14]
  wire  geu; // @[BrCond.scala 44:14]
  wire  _T_7; // @[BrCond.scala 46:18]
  wire  _T_8; // @[BrCond.scala 46:29]
  wire  _T_9; // @[BrCond.scala 47:18]
  wire  _T_10; // @[BrCond.scala 47:29]
  wire  _T_11; // @[BrCond.scala 46:36]
  wire  _T_12; // @[BrCond.scala 48:18]
  wire  _T_13; // @[BrCond.scala 48:29]
  wire  _T_14; // @[BrCond.scala 47:37]
  wire  _T_15; // @[BrCond.scala 49:18]
  wire  _T_16; // @[BrCond.scala 49:29]
  wire  _T_17; // @[BrCond.scala 48:36]
  wire  _T_18; // @[BrCond.scala 50:18]
  wire  _T_19; // @[BrCond.scala 50:30]
  wire  _T_20; // @[BrCond.scala 49:36]
  wire  _T_21; // @[BrCond.scala 51:18]
  wire  _T_22; // @[BrCond.scala 51:30]
  assign diff = io_rs1 - io_rs2; // @[BrCond.scala 37:21]
  assign neq = diff != 32'h0; // @[BrCond.scala 38:19]
  assign eq = neq == 1'h0; // @[BrCond.scala 39:14]
  assign _T_1 = io_rs1[31]; // @[BrCond.scala 40:26]
  assign _T_2 = io_rs2[31]; // @[BrCond.scala 40:45]
  assign isSameSign = _T_1 == _T_2; // @[BrCond.scala 40:35]
  assign _T_3 = diff[31]; // @[BrCond.scala 41:34]
  assign lt = isSameSign ? _T_3 : _T_1; // @[BrCond.scala 41:17]
  assign ltu = isSameSign ? _T_3 : _T_2; // @[BrCond.scala 42:17]
  assign ge = lt == 1'h0; // @[BrCond.scala 43:14]
  assign geu = ltu == 1'h0; // @[BrCond.scala 44:14]
  assign _T_7 = io_br_type == 3'h3; // @[BrCond.scala 46:18]
  assign _T_8 = _T_7 & eq; // @[BrCond.scala 46:29]
  assign _T_9 = io_br_type == 3'h6; // @[BrCond.scala 47:18]
  assign _T_10 = _T_9 & neq; // @[BrCond.scala 47:29]
  assign _T_11 = _T_8 | _T_10; // @[BrCond.scala 46:36]
  assign _T_12 = io_br_type == 3'h2; // @[BrCond.scala 48:18]
  assign _T_13 = _T_12 & lt; // @[BrCond.scala 48:29]
  assign _T_14 = _T_11 | _T_13; // @[BrCond.scala 47:37]
  assign _T_15 = io_br_type == 3'h5; // @[BrCond.scala 49:18]
  assign _T_16 = _T_15 & ge; // @[BrCond.scala 49:29]
  assign _T_17 = _T_14 | _T_16; // @[BrCond.scala 48:36]
  assign _T_18 = io_br_type == 3'h1; // @[BrCond.scala 50:18]
  assign _T_19 = _T_18 & ltu; // @[BrCond.scala 50:30]
  assign _T_20 = _T_17 | _T_19; // @[BrCond.scala 49:36]
  assign _T_21 = io_br_type == 3'h4; // @[BrCond.scala 51:18]
  assign _T_22 = _T_21 & geu; // @[BrCond.scala 51:30]
  assign io_taken = _T_20 | _T_22; // @[BrCond.scala 45:12]
endmodule
