module ImmGenWire(
  input  [31:0] io_inst,
  input  [2:0]  io_sel,
  output [31:0] io_out
);
  wire [11:0] _T; // @[ImmGen.scala 21:21]
  wire [11:0] Iimm; // @[ImmGen.scala 21:30]
  wire [6:0] _T_1; // @[ImmGen.scala 22:25]
  wire [4:0] _T_2; // @[ImmGen.scala 22:42]
  wire [11:0] _T_3; // @[Cat.scala 29:58]
  wire [11:0] Simm; // @[ImmGen.scala 22:50]
  wire  _T_4; // @[ImmGen.scala 23:25]
  wire  _T_5; // @[ImmGen.scala 23:38]
  wire [5:0] _T_6; // @[ImmGen.scala 23:50]
  wire [3:0] _T_7; // @[ImmGen.scala 23:67]
  wire [12:0] _T_11; // @[Cat.scala 29:58]
  wire [12:0] Bimm; // @[ImmGen.scala 23:86]
  wire [19:0] _T_12; // @[ImmGen.scala 24:25]
  wire [31:0] _T_13; // @[Cat.scala 29:58]
  wire [31:0] Uimm; // @[ImmGen.scala 24:46]
  wire [7:0] _T_15; // @[ImmGen.scala 25:38]
  wire  _T_16; // @[ImmGen.scala 25:55]
  wire [3:0] _T_18; // @[ImmGen.scala 25:85]
  wire [20:0] _T_23; // @[Cat.scala 29:58]
  wire [20:0] Jimm; // @[ImmGen.scala 25:105]
  wire [4:0] _T_24; // @[ImmGen.scala 26:21]
  wire [5:0] Zimm; // @[ImmGen.scala 26:30]
  wire [11:0] _T_25; // @[ImmGen.scala 28:36]
  wire [11:0] _T_26; // @[ImmGen.scala 28:36]
  wire  _T_27; // @[Mux.scala 80:60]
  wire [11:0] _T_28; // @[Mux.scala 80:57]
  wire  _T_29; // @[Mux.scala 80:60]
  wire [11:0] _T_30; // @[Mux.scala 80:57]
  wire  _T_31; // @[Mux.scala 80:60]
  wire [12:0] _T_32; // @[Mux.scala 80:57]
  wire  _T_33; // @[Mux.scala 80:60]
  wire [31:0] _T_34; // @[Mux.scala 80:57]
  wire  _T_35; // @[Mux.scala 80:60]
  wire [31:0] _T_36; // @[Mux.scala 80:57]
  wire  _T_37; // @[Mux.scala 80:60]
  wire [31:0] _T_38; // @[Mux.scala 80:57]
  assign _T = io_inst[31:20]; // @[ImmGen.scala 21:21]
  assign Iimm = $signed(_T); // @[ImmGen.scala 21:30]
  assign _T_1 = io_inst[31:25]; // @[ImmGen.scala 22:25]
  assign _T_2 = io_inst[11:7]; // @[ImmGen.scala 22:42]
  assign _T_3 = {_T_1,_T_2}; // @[Cat.scala 29:58]
  assign Simm = $signed(_T_3); // @[ImmGen.scala 22:50]
  assign _T_4 = io_inst[31]; // @[ImmGen.scala 23:25]
  assign _T_5 = io_inst[7]; // @[ImmGen.scala 23:38]
  assign _T_6 = io_inst[30:25]; // @[ImmGen.scala 23:50]
  assign _T_7 = io_inst[11:8]; // @[ImmGen.scala 23:67]
  assign _T_11 = {_T_4,_T_5,_T_6,_T_7,1'h0}; // @[Cat.scala 29:58]
  assign Bimm = $signed(_T_11); // @[ImmGen.scala 23:86]
  assign _T_12 = io_inst[31:12]; // @[ImmGen.scala 24:25]
  assign _T_13 = {_T_12,12'h0}; // @[Cat.scala 29:58]
  assign Uimm = $signed(_T_13); // @[ImmGen.scala 24:46]
  assign _T_15 = io_inst[19:12]; // @[ImmGen.scala 25:38]
  assign _T_16 = io_inst[20]; // @[ImmGen.scala 25:55]
  assign _T_18 = io_inst[24:21]; // @[ImmGen.scala 25:85]
  assign _T_23 = {_T_4,_T_15,_T_16,_T_6,_T_18,1'h0}; // @[Cat.scala 29:58]
  assign Jimm = $signed(_T_23); // @[ImmGen.scala 25:105]
  assign _T_24 = io_inst[19:15]; // @[ImmGen.scala 26:21]
  assign Zimm = {1'b0,$signed(_T_24)}; // @[ImmGen.scala 26:30]
  assign _T_25 = $signed(Iimm) & $signed(-12'sh2); // @[ImmGen.scala 28:36]
  assign _T_26 = $signed(_T_25); // @[ImmGen.scala 28:36]
  assign _T_27 = 3'h1 == io_sel; // @[Mux.scala 80:60]
  assign _T_28 = _T_27 ? $signed(Iimm) : $signed(_T_26); // @[Mux.scala 80:57]
  assign _T_29 = 3'h2 == io_sel; // @[Mux.scala 80:60]
  assign _T_30 = _T_29 ? $signed(Simm) : $signed(_T_28); // @[Mux.scala 80:57]
  assign _T_31 = 3'h5 == io_sel; // @[Mux.scala 80:60]
  assign _T_32 = _T_31 ? $signed(Bimm) : $signed({{1{_T_30[11]}},_T_30}); // @[Mux.scala 80:57]
  assign _T_33 = 3'h3 == io_sel; // @[Mux.scala 80:60]
  assign _T_34 = _T_33 ? $signed(Uimm) : $signed({{19{_T_32[12]}},_T_32}); // @[Mux.scala 80:57]
  assign _T_35 = 3'h4 == io_sel; // @[Mux.scala 80:60]
  assign _T_36 = _T_35 ? $signed({{11{Jimm[20]}},Jimm}) : $signed(_T_34); // @[Mux.scala 80:57]
  assign _T_37 = 3'h6 == io_sel; // @[Mux.scala 80:60]
  assign _T_38 = _T_37 ? $signed({{26{Zimm[5]}},Zimm}) : $signed(_T_36); // @[Mux.scala 80:57]
  assign io_out = $unsigned(_T_38); // @[ImmGen.scala 28:10]
endmodule
