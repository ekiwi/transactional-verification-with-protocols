module Control(
  input  [31:0] io_inst,
  output [1:0]  io_pc_sel,
  output        io_inst_kill,
  output        io_A_sel,
  output        io_B_sel,
  output [2:0]  io_imm_sel,
  output [3:0]  io_alu_op,
  output [2:0]  io_br_type,
  output [1:0]  io_st_type,
  output [2:0]  io_ld_type,
  output [1:0]  io_wb_sel,
  output        io_wb_en,
  output [2:0]  io_csr_cmd,
  output        io_illegal
);
  wire [31:0] _T; // @[Lookup.scala 31:38]
  wire  _T_1; // @[Lookup.scala 31:38]
  wire  _T_3; // @[Lookup.scala 31:38]
  wire  _T_5; // @[Lookup.scala 31:38]
  wire [31:0] _T_6; // @[Lookup.scala 31:38]
  wire  _T_7; // @[Lookup.scala 31:38]
  wire  _T_9; // @[Lookup.scala 31:38]
  wire  _T_11; // @[Lookup.scala 31:38]
  wire  _T_13; // @[Lookup.scala 31:38]
  wire  _T_15; // @[Lookup.scala 31:38]
  wire  _T_17; // @[Lookup.scala 31:38]
  wire  _T_19; // @[Lookup.scala 31:38]
  wire  _T_21; // @[Lookup.scala 31:38]
  wire  _T_23; // @[Lookup.scala 31:38]
  wire  _T_25; // @[Lookup.scala 31:38]
  wire  _T_27; // @[Lookup.scala 31:38]
  wire  _T_29; // @[Lookup.scala 31:38]
  wire  _T_31; // @[Lookup.scala 31:38]
  wire  _T_33; // @[Lookup.scala 31:38]
  wire  _T_35; // @[Lookup.scala 31:38]
  wire  _T_37; // @[Lookup.scala 31:38]
  wire  _T_39; // @[Lookup.scala 31:38]
  wire  _T_41; // @[Lookup.scala 31:38]
  wire  _T_43; // @[Lookup.scala 31:38]
  wire  _T_45; // @[Lookup.scala 31:38]
  wire  _T_47; // @[Lookup.scala 31:38]
  wire [31:0] _T_48; // @[Lookup.scala 31:38]
  wire  _T_49; // @[Lookup.scala 31:38]
  wire  _T_51; // @[Lookup.scala 31:38]
  wire  _T_53; // @[Lookup.scala 31:38]
  wire  _T_55; // @[Lookup.scala 31:38]
  wire  _T_57; // @[Lookup.scala 31:38]
  wire  _T_59; // @[Lookup.scala 31:38]
  wire  _T_61; // @[Lookup.scala 31:38]
  wire  _T_63; // @[Lookup.scala 31:38]
  wire  _T_65; // @[Lookup.scala 31:38]
  wire  _T_67; // @[Lookup.scala 31:38]
  wire  _T_69; // @[Lookup.scala 31:38]
  wire  _T_71; // @[Lookup.scala 31:38]
  wire  _T_73; // @[Lookup.scala 31:38]
  wire [31:0] _T_74; // @[Lookup.scala 31:38]
  wire  _T_75; // @[Lookup.scala 31:38]
  wire  _T_77; // @[Lookup.scala 31:38]
  wire  _T_79; // @[Lookup.scala 31:38]
  wire  _T_81; // @[Lookup.scala 31:38]
  wire  _T_83; // @[Lookup.scala 31:38]
  wire  _T_85; // @[Lookup.scala 31:38]
  wire  _T_87; // @[Lookup.scala 31:38]
  wire  _T_89; // @[Lookup.scala 31:38]
  wire  _T_91; // @[Lookup.scala 31:38]
  wire  _T_93; // @[Lookup.scala 31:38]
  wire  _T_95; // @[Lookup.scala 31:38]
  wire  _T_97; // @[Lookup.scala 31:38]
  wire [1:0] _T_99; // @[Lookup.scala 33:37]
  wire [1:0] _T_100; // @[Lookup.scala 33:37]
  wire [1:0] _T_101; // @[Lookup.scala 33:37]
  wire [1:0] _T_102; // @[Lookup.scala 33:37]
  wire [1:0] _T_103; // @[Lookup.scala 33:37]
  wire [1:0] _T_104; // @[Lookup.scala 33:37]
  wire [1:0] _T_105; // @[Lookup.scala 33:37]
  wire [1:0] _T_106; // @[Lookup.scala 33:37]
  wire [1:0] _T_107; // @[Lookup.scala 33:37]
  wire [1:0] _T_108; // @[Lookup.scala 33:37]
  wire [1:0] _T_109; // @[Lookup.scala 33:37]
  wire [1:0] _T_110; // @[Lookup.scala 33:37]
  wire [1:0] _T_111; // @[Lookup.scala 33:37]
  wire [1:0] _T_112; // @[Lookup.scala 33:37]
  wire [1:0] _T_113; // @[Lookup.scala 33:37]
  wire [1:0] _T_114; // @[Lookup.scala 33:37]
  wire [1:0] _T_115; // @[Lookup.scala 33:37]
  wire [1:0] _T_116; // @[Lookup.scala 33:37]
  wire [1:0] _T_117; // @[Lookup.scala 33:37]
  wire [1:0] _T_118; // @[Lookup.scala 33:37]
  wire [1:0] _T_119; // @[Lookup.scala 33:37]
  wire [1:0] _T_120; // @[Lookup.scala 33:37]
  wire [1:0] _T_121; // @[Lookup.scala 33:37]
  wire [1:0] _T_122; // @[Lookup.scala 33:37]
  wire [1:0] _T_123; // @[Lookup.scala 33:37]
  wire [1:0] _T_124; // @[Lookup.scala 33:37]
  wire [1:0] _T_125; // @[Lookup.scala 33:37]
  wire [1:0] _T_126; // @[Lookup.scala 33:37]
  wire [1:0] _T_127; // @[Lookup.scala 33:37]
  wire [1:0] _T_128; // @[Lookup.scala 33:37]
  wire [1:0] _T_129; // @[Lookup.scala 33:37]
  wire [1:0] _T_130; // @[Lookup.scala 33:37]
  wire [1:0] _T_131; // @[Lookup.scala 33:37]
  wire [1:0] _T_132; // @[Lookup.scala 33:37]
  wire [1:0] _T_133; // @[Lookup.scala 33:37]
  wire [1:0] _T_134; // @[Lookup.scala 33:37]
  wire [1:0] _T_135; // @[Lookup.scala 33:37]
  wire [1:0] _T_136; // @[Lookup.scala 33:37]
  wire [1:0] _T_137; // @[Lookup.scala 33:37]
  wire [1:0] _T_138; // @[Lookup.scala 33:37]
  wire [1:0] _T_139; // @[Lookup.scala 33:37]
  wire [1:0] _T_140; // @[Lookup.scala 33:37]
  wire [1:0] _T_141; // @[Lookup.scala 33:37]
  wire [1:0] _T_142; // @[Lookup.scala 33:37]
  wire [1:0] _T_143; // @[Lookup.scala 33:37]
  wire [1:0] _T_144; // @[Lookup.scala 33:37]
  wire [1:0] _T_145; // @[Lookup.scala 33:37]
  wire  _T_154; // @[Lookup.scala 33:37]
  wire  _T_155; // @[Lookup.scala 33:37]
  wire  _T_156; // @[Lookup.scala 33:37]
  wire  _T_157; // @[Lookup.scala 33:37]
  wire  _T_158; // @[Lookup.scala 33:37]
  wire  _T_159; // @[Lookup.scala 33:37]
  wire  _T_160; // @[Lookup.scala 33:37]
  wire  _T_161; // @[Lookup.scala 33:37]
  wire  _T_162; // @[Lookup.scala 33:37]
  wire  _T_163; // @[Lookup.scala 33:37]
  wire  _T_164; // @[Lookup.scala 33:37]
  wire  _T_165; // @[Lookup.scala 33:37]
  wire  _T_166; // @[Lookup.scala 33:37]
  wire  _T_167; // @[Lookup.scala 33:37]
  wire  _T_168; // @[Lookup.scala 33:37]
  wire  _T_169; // @[Lookup.scala 33:37]
  wire  _T_170; // @[Lookup.scala 33:37]
  wire  _T_171; // @[Lookup.scala 33:37]
  wire  _T_172; // @[Lookup.scala 33:37]
  wire  _T_173; // @[Lookup.scala 33:37]
  wire  _T_174; // @[Lookup.scala 33:37]
  wire  _T_175; // @[Lookup.scala 33:37]
  wire  _T_176; // @[Lookup.scala 33:37]
  wire  _T_177; // @[Lookup.scala 33:37]
  wire  _T_178; // @[Lookup.scala 33:37]
  wire  _T_179; // @[Lookup.scala 33:37]
  wire  _T_180; // @[Lookup.scala 33:37]
  wire  _T_181; // @[Lookup.scala 33:37]
  wire  _T_182; // @[Lookup.scala 33:37]
  wire  _T_183; // @[Lookup.scala 33:37]
  wire  _T_184; // @[Lookup.scala 33:37]
  wire  _T_185; // @[Lookup.scala 33:37]
  wire  _T_186; // @[Lookup.scala 33:37]
  wire  _T_187; // @[Lookup.scala 33:37]
  wire  _T_188; // @[Lookup.scala 33:37]
  wire  _T_189; // @[Lookup.scala 33:37]
  wire  _T_190; // @[Lookup.scala 33:37]
  wire  _T_191; // @[Lookup.scala 33:37]
  wire  _T_192; // @[Lookup.scala 33:37]
  wire  _T_193; // @[Lookup.scala 33:37]
  wire  _T_207; // @[Lookup.scala 33:37]
  wire  _T_208; // @[Lookup.scala 33:37]
  wire  _T_209; // @[Lookup.scala 33:37]
  wire  _T_210; // @[Lookup.scala 33:37]
  wire  _T_211; // @[Lookup.scala 33:37]
  wire  _T_212; // @[Lookup.scala 33:37]
  wire  _T_213; // @[Lookup.scala 33:37]
  wire  _T_214; // @[Lookup.scala 33:37]
  wire  _T_215; // @[Lookup.scala 33:37]
  wire  _T_216; // @[Lookup.scala 33:37]
  wire  _T_217; // @[Lookup.scala 33:37]
  wire  _T_218; // @[Lookup.scala 33:37]
  wire  _T_219; // @[Lookup.scala 33:37]
  wire  _T_220; // @[Lookup.scala 33:37]
  wire  _T_221; // @[Lookup.scala 33:37]
  wire  _T_222; // @[Lookup.scala 33:37]
  wire  _T_223; // @[Lookup.scala 33:37]
  wire  _T_224; // @[Lookup.scala 33:37]
  wire  _T_225; // @[Lookup.scala 33:37]
  wire  _T_226; // @[Lookup.scala 33:37]
  wire  _T_227; // @[Lookup.scala 33:37]
  wire  _T_228; // @[Lookup.scala 33:37]
  wire  _T_229; // @[Lookup.scala 33:37]
  wire  _T_230; // @[Lookup.scala 33:37]
  wire  _T_231; // @[Lookup.scala 33:37]
  wire  _T_232; // @[Lookup.scala 33:37]
  wire  _T_233; // @[Lookup.scala 33:37]
  wire  _T_234; // @[Lookup.scala 33:37]
  wire  _T_235; // @[Lookup.scala 33:37]
  wire  _T_236; // @[Lookup.scala 33:37]
  wire  _T_237; // @[Lookup.scala 33:37]
  wire  _T_238; // @[Lookup.scala 33:37]
  wire  _T_239; // @[Lookup.scala 33:37]
  wire  _T_240; // @[Lookup.scala 33:37]
  wire  _T_241; // @[Lookup.scala 33:37]
  wire [2:0] _T_246; // @[Lookup.scala 33:37]
  wire [2:0] _T_247; // @[Lookup.scala 33:37]
  wire [2:0] _T_248; // @[Lookup.scala 33:37]
  wire [2:0] _T_249; // @[Lookup.scala 33:37]
  wire [2:0] _T_250; // @[Lookup.scala 33:37]
  wire [2:0] _T_251; // @[Lookup.scala 33:37]
  wire [2:0] _T_252; // @[Lookup.scala 33:37]
  wire [2:0] _T_253; // @[Lookup.scala 33:37]
  wire [2:0] _T_254; // @[Lookup.scala 33:37]
  wire [2:0] _T_255; // @[Lookup.scala 33:37]
  wire [2:0] _T_256; // @[Lookup.scala 33:37]
  wire [2:0] _T_257; // @[Lookup.scala 33:37]
  wire [2:0] _T_258; // @[Lookup.scala 33:37]
  wire [2:0] _T_259; // @[Lookup.scala 33:37]
  wire [2:0] _T_260; // @[Lookup.scala 33:37]
  wire [2:0] _T_261; // @[Lookup.scala 33:37]
  wire [2:0] _T_262; // @[Lookup.scala 33:37]
  wire [2:0] _T_263; // @[Lookup.scala 33:37]
  wire [2:0] _T_264; // @[Lookup.scala 33:37]
  wire [2:0] _T_265; // @[Lookup.scala 33:37]
  wire [2:0] _T_266; // @[Lookup.scala 33:37]
  wire [2:0] _T_267; // @[Lookup.scala 33:37]
  wire [2:0] _T_268; // @[Lookup.scala 33:37]
  wire [2:0] _T_269; // @[Lookup.scala 33:37]
  wire [2:0] _T_270; // @[Lookup.scala 33:37]
  wire [2:0] _T_271; // @[Lookup.scala 33:37]
  wire [2:0] _T_272; // @[Lookup.scala 33:37]
  wire [2:0] _T_273; // @[Lookup.scala 33:37]
  wire [2:0] _T_274; // @[Lookup.scala 33:37]
  wire [2:0] _T_275; // @[Lookup.scala 33:37]
  wire [2:0] _T_276; // @[Lookup.scala 33:37]
  wire [2:0] _T_277; // @[Lookup.scala 33:37]
  wire [2:0] _T_278; // @[Lookup.scala 33:37]
  wire [2:0] _T_279; // @[Lookup.scala 33:37]
  wire [2:0] _T_280; // @[Lookup.scala 33:37]
  wire [2:0] _T_281; // @[Lookup.scala 33:37]
  wire [2:0] _T_282; // @[Lookup.scala 33:37]
  wire [2:0] _T_283; // @[Lookup.scala 33:37]
  wire [2:0] _T_284; // @[Lookup.scala 33:37]
  wire [2:0] _T_285; // @[Lookup.scala 33:37]
  wire [2:0] _T_286; // @[Lookup.scala 33:37]
  wire [2:0] _T_287; // @[Lookup.scala 33:37]
  wire [2:0] _T_288; // @[Lookup.scala 33:37]
  wire [2:0] _T_289; // @[Lookup.scala 33:37]
  wire [3:0] _T_297; // @[Lookup.scala 33:37]
  wire [3:0] _T_298; // @[Lookup.scala 33:37]
  wire [3:0] _T_299; // @[Lookup.scala 33:37]
  wire [3:0] _T_300; // @[Lookup.scala 33:37]
  wire [3:0] _T_301; // @[Lookup.scala 33:37]
  wire [3:0] _T_302; // @[Lookup.scala 33:37]
  wire [3:0] _T_303; // @[Lookup.scala 33:37]
  wire [3:0] _T_304; // @[Lookup.scala 33:37]
  wire [3:0] _T_305; // @[Lookup.scala 33:37]
  wire [3:0] _T_306; // @[Lookup.scala 33:37]
  wire [3:0] _T_307; // @[Lookup.scala 33:37]
  wire [3:0] _T_308; // @[Lookup.scala 33:37]
  wire [3:0] _T_309; // @[Lookup.scala 33:37]
  wire [3:0] _T_310; // @[Lookup.scala 33:37]
  wire [3:0] _T_311; // @[Lookup.scala 33:37]
  wire [3:0] _T_312; // @[Lookup.scala 33:37]
  wire [3:0] _T_313; // @[Lookup.scala 33:37]
  wire [3:0] _T_314; // @[Lookup.scala 33:37]
  wire [3:0] _T_315; // @[Lookup.scala 33:37]
  wire [3:0] _T_316; // @[Lookup.scala 33:37]
  wire [3:0] _T_317; // @[Lookup.scala 33:37]
  wire [3:0] _T_318; // @[Lookup.scala 33:37]
  wire [3:0] _T_319; // @[Lookup.scala 33:37]
  wire [3:0] _T_320; // @[Lookup.scala 33:37]
  wire [3:0] _T_321; // @[Lookup.scala 33:37]
  wire [3:0] _T_322; // @[Lookup.scala 33:37]
  wire [3:0] _T_323; // @[Lookup.scala 33:37]
  wire [3:0] _T_324; // @[Lookup.scala 33:37]
  wire [3:0] _T_325; // @[Lookup.scala 33:37]
  wire [3:0] _T_326; // @[Lookup.scala 33:37]
  wire [3:0] _T_327; // @[Lookup.scala 33:37]
  wire [3:0] _T_328; // @[Lookup.scala 33:37]
  wire [3:0] _T_329; // @[Lookup.scala 33:37]
  wire [3:0] _T_330; // @[Lookup.scala 33:37]
  wire [3:0] _T_331; // @[Lookup.scala 33:37]
  wire [3:0] _T_332; // @[Lookup.scala 33:37]
  wire [3:0] _T_333; // @[Lookup.scala 33:37]
  wire [3:0] _T_334; // @[Lookup.scala 33:37]
  wire [3:0] _T_335; // @[Lookup.scala 33:37]
  wire [3:0] _T_336; // @[Lookup.scala 33:37]
  wire [3:0] _T_337; // @[Lookup.scala 33:37]
  wire [2:0] _T_377; // @[Lookup.scala 33:37]
  wire [2:0] _T_378; // @[Lookup.scala 33:37]
  wire [2:0] _T_379; // @[Lookup.scala 33:37]
  wire [2:0] _T_380; // @[Lookup.scala 33:37]
  wire [2:0] _T_381; // @[Lookup.scala 33:37]
  wire [2:0] _T_382; // @[Lookup.scala 33:37]
  wire [2:0] _T_383; // @[Lookup.scala 33:37]
  wire [2:0] _T_384; // @[Lookup.scala 33:37]
  wire [2:0] _T_385; // @[Lookup.scala 33:37]
  wire  _T_388; // @[Lookup.scala 33:37]
  wire  _T_389; // @[Lookup.scala 33:37]
  wire  _T_390; // @[Lookup.scala 33:37]
  wire  _T_391; // @[Lookup.scala 33:37]
  wire  _T_392; // @[Lookup.scala 33:37]
  wire  _T_393; // @[Lookup.scala 33:37]
  wire  _T_394; // @[Lookup.scala 33:37]
  wire  _T_395; // @[Lookup.scala 33:37]
  wire  _T_396; // @[Lookup.scala 33:37]
  wire  _T_397; // @[Lookup.scala 33:37]
  wire  _T_398; // @[Lookup.scala 33:37]
  wire  _T_399; // @[Lookup.scala 33:37]
  wire  _T_400; // @[Lookup.scala 33:37]
  wire  _T_401; // @[Lookup.scala 33:37]
  wire  _T_402; // @[Lookup.scala 33:37]
  wire  _T_403; // @[Lookup.scala 33:37]
  wire  _T_404; // @[Lookup.scala 33:37]
  wire  _T_405; // @[Lookup.scala 33:37]
  wire  _T_406; // @[Lookup.scala 33:37]
  wire  _T_407; // @[Lookup.scala 33:37]
  wire  _T_408; // @[Lookup.scala 33:37]
  wire  _T_409; // @[Lookup.scala 33:37]
  wire  _T_410; // @[Lookup.scala 33:37]
  wire  _T_411; // @[Lookup.scala 33:37]
  wire  _T_412; // @[Lookup.scala 33:37]
  wire  _T_413; // @[Lookup.scala 33:37]
  wire  _T_414; // @[Lookup.scala 33:37]
  wire  _T_415; // @[Lookup.scala 33:37]
  wire  _T_416; // @[Lookup.scala 33:37]
  wire  _T_417; // @[Lookup.scala 33:37]
  wire  _T_418; // @[Lookup.scala 33:37]
  wire  _T_419; // @[Lookup.scala 33:37]
  wire  _T_420; // @[Lookup.scala 33:37]
  wire  _T_421; // @[Lookup.scala 33:37]
  wire  _T_422; // @[Lookup.scala 33:37]
  wire  _T_423; // @[Lookup.scala 33:37]
  wire  _T_424; // @[Lookup.scala 33:37]
  wire  _T_425; // @[Lookup.scala 33:37]
  wire  _T_426; // @[Lookup.scala 33:37]
  wire  _T_427; // @[Lookup.scala 33:37]
  wire  _T_428; // @[Lookup.scala 33:37]
  wire  _T_429; // @[Lookup.scala 33:37]
  wire  _T_430; // @[Lookup.scala 33:37]
  wire  _T_431; // @[Lookup.scala 33:37]
  wire  _T_432; // @[Lookup.scala 33:37]
  wire  _T_433; // @[Lookup.scala 33:37]
  wire [1:0] _T_465; // @[Lookup.scala 33:37]
  wire [1:0] _T_466; // @[Lookup.scala 33:37]
  wire [1:0] _T_467; // @[Lookup.scala 33:37]
  wire [1:0] _T_468; // @[Lookup.scala 33:37]
  wire [1:0] _T_469; // @[Lookup.scala 33:37]
  wire [1:0] _T_470; // @[Lookup.scala 33:37]
  wire [1:0] _T_471; // @[Lookup.scala 33:37]
  wire [1:0] _T_472; // @[Lookup.scala 33:37]
  wire [1:0] _T_473; // @[Lookup.scala 33:37]
  wire [1:0] _T_474; // @[Lookup.scala 33:37]
  wire [1:0] _T_475; // @[Lookup.scala 33:37]
  wire [1:0] _T_476; // @[Lookup.scala 33:37]
  wire [1:0] _T_477; // @[Lookup.scala 33:37]
  wire [1:0] _T_478; // @[Lookup.scala 33:37]
  wire [1:0] _T_479; // @[Lookup.scala 33:37]
  wire [1:0] _T_480; // @[Lookup.scala 33:37]
  wire [1:0] _T_481; // @[Lookup.scala 33:37]
  wire [2:0] _T_516; // @[Lookup.scala 33:37]
  wire [2:0] _T_517; // @[Lookup.scala 33:37]
  wire [2:0] _T_518; // @[Lookup.scala 33:37]
  wire [2:0] _T_519; // @[Lookup.scala 33:37]
  wire [2:0] _T_520; // @[Lookup.scala 33:37]
  wire [2:0] _T_521; // @[Lookup.scala 33:37]
  wire [2:0] _T_522; // @[Lookup.scala 33:37]
  wire [2:0] _T_523; // @[Lookup.scala 33:37]
  wire [2:0] _T_524; // @[Lookup.scala 33:37]
  wire [2:0] _T_525; // @[Lookup.scala 33:37]
  wire [2:0] _T_526; // @[Lookup.scala 33:37]
  wire [2:0] _T_527; // @[Lookup.scala 33:37]
  wire [2:0] _T_528; // @[Lookup.scala 33:37]
  wire [2:0] _T_529; // @[Lookup.scala 33:37]
  wire [1:0] _T_532; // @[Lookup.scala 33:37]
  wire [1:0] _T_533; // @[Lookup.scala 33:37]
  wire [1:0] _T_534; // @[Lookup.scala 33:37]
  wire [1:0] _T_535; // @[Lookup.scala 33:37]
  wire [1:0] _T_536; // @[Lookup.scala 33:37]
  wire [1:0] _T_537; // @[Lookup.scala 33:37]
  wire [1:0] _T_538; // @[Lookup.scala 33:37]
  wire [1:0] _T_539; // @[Lookup.scala 33:37]
  wire [1:0] _T_540; // @[Lookup.scala 33:37]
  wire [1:0] _T_541; // @[Lookup.scala 33:37]
  wire [1:0] _T_542; // @[Lookup.scala 33:37]
  wire [1:0] _T_543; // @[Lookup.scala 33:37]
  wire [1:0] _T_544; // @[Lookup.scala 33:37]
  wire [1:0] _T_545; // @[Lookup.scala 33:37]
  wire [1:0] _T_546; // @[Lookup.scala 33:37]
  wire [1:0] _T_547; // @[Lookup.scala 33:37]
  wire [1:0] _T_548; // @[Lookup.scala 33:37]
  wire [1:0] _T_549; // @[Lookup.scala 33:37]
  wire [1:0] _T_550; // @[Lookup.scala 33:37]
  wire [1:0] _T_551; // @[Lookup.scala 33:37]
  wire [1:0] _T_552; // @[Lookup.scala 33:37]
  wire [1:0] _T_553; // @[Lookup.scala 33:37]
  wire [1:0] _T_554; // @[Lookup.scala 33:37]
  wire [1:0] _T_555; // @[Lookup.scala 33:37]
  wire [1:0] _T_556; // @[Lookup.scala 33:37]
  wire [1:0] _T_557; // @[Lookup.scala 33:37]
  wire [1:0] _T_558; // @[Lookup.scala 33:37]
  wire [1:0] _T_559; // @[Lookup.scala 33:37]
  wire [1:0] _T_560; // @[Lookup.scala 33:37]
  wire [1:0] _T_561; // @[Lookup.scala 33:37]
  wire [1:0] _T_562; // @[Lookup.scala 33:37]
  wire [1:0] _T_563; // @[Lookup.scala 33:37]
  wire [1:0] _T_564; // @[Lookup.scala 33:37]
  wire [1:0] _T_565; // @[Lookup.scala 33:37]
  wire [1:0] _T_566; // @[Lookup.scala 33:37]
  wire [1:0] _T_567; // @[Lookup.scala 33:37]
  wire [1:0] _T_568; // @[Lookup.scala 33:37]
  wire [1:0] _T_569; // @[Lookup.scala 33:37]
  wire [1:0] _T_570; // @[Lookup.scala 33:37]
  wire [1:0] _T_571; // @[Lookup.scala 33:37]
  wire [1:0] _T_572; // @[Lookup.scala 33:37]
  wire [1:0] _T_573; // @[Lookup.scala 33:37]
  wire [1:0] _T_574; // @[Lookup.scala 33:37]
  wire [1:0] _T_575; // @[Lookup.scala 33:37]
  wire [1:0] _T_576; // @[Lookup.scala 33:37]
  wire [1:0] _T_577; // @[Lookup.scala 33:37]
  wire  _T_583; // @[Lookup.scala 33:37]
  wire  _T_584; // @[Lookup.scala 33:37]
  wire  _T_585; // @[Lookup.scala 33:37]
  wire  _T_586; // @[Lookup.scala 33:37]
  wire  _T_587; // @[Lookup.scala 33:37]
  wire  _T_588; // @[Lookup.scala 33:37]
  wire  _T_589; // @[Lookup.scala 33:37]
  wire  _T_590; // @[Lookup.scala 33:37]
  wire  _T_591; // @[Lookup.scala 33:37]
  wire  _T_592; // @[Lookup.scala 33:37]
  wire  _T_593; // @[Lookup.scala 33:37]
  wire  _T_594; // @[Lookup.scala 33:37]
  wire  _T_595; // @[Lookup.scala 33:37]
  wire  _T_596; // @[Lookup.scala 33:37]
  wire  _T_597; // @[Lookup.scala 33:37]
  wire  _T_598; // @[Lookup.scala 33:37]
  wire  _T_599; // @[Lookup.scala 33:37]
  wire  _T_600; // @[Lookup.scala 33:37]
  wire  _T_601; // @[Lookup.scala 33:37]
  wire  _T_602; // @[Lookup.scala 33:37]
  wire  _T_603; // @[Lookup.scala 33:37]
  wire  _T_604; // @[Lookup.scala 33:37]
  wire  _T_605; // @[Lookup.scala 33:37]
  wire  _T_606; // @[Lookup.scala 33:37]
  wire  _T_607; // @[Lookup.scala 33:37]
  wire  _T_608; // @[Lookup.scala 33:37]
  wire  _T_609; // @[Lookup.scala 33:37]
  wire  _T_610; // @[Lookup.scala 33:37]
  wire  _T_611; // @[Lookup.scala 33:37]
  wire  _T_612; // @[Lookup.scala 33:37]
  wire  _T_613; // @[Lookup.scala 33:37]
  wire  _T_614; // @[Lookup.scala 33:37]
  wire  _T_615; // @[Lookup.scala 33:37]
  wire  _T_616; // @[Lookup.scala 33:37]
  wire  _T_617; // @[Lookup.scala 33:37]
  wire  _T_618; // @[Lookup.scala 33:37]
  wire  _T_619; // @[Lookup.scala 33:37]
  wire  _T_620; // @[Lookup.scala 33:37]
  wire  _T_621; // @[Lookup.scala 33:37]
  wire  _T_622; // @[Lookup.scala 33:37]
  wire  _T_623; // @[Lookup.scala 33:37]
  wire  _T_624; // @[Lookup.scala 33:37]
  wire  _T_625; // @[Lookup.scala 33:37]
  wire [2:0] _T_627; // @[Lookup.scala 33:37]
  wire [2:0] _T_628; // @[Lookup.scala 33:37]
  wire [2:0] _T_629; // @[Lookup.scala 33:37]
  wire [2:0] _T_630; // @[Lookup.scala 33:37]
  wire [2:0] _T_631; // @[Lookup.scala 33:37]
  wire [2:0] _T_632; // @[Lookup.scala 33:37]
  wire [2:0] _T_633; // @[Lookup.scala 33:37]
  wire [2:0] _T_634; // @[Lookup.scala 33:37]
  wire [2:0] _T_635; // @[Lookup.scala 33:37]
  wire [2:0] _T_636; // @[Lookup.scala 33:37]
  wire [2:0] _T_637; // @[Lookup.scala 33:37]
  wire [2:0] _T_638; // @[Lookup.scala 33:37]
  wire [2:0] _T_639; // @[Lookup.scala 33:37]
  wire [2:0] _T_640; // @[Lookup.scala 33:37]
  wire [2:0] _T_641; // @[Lookup.scala 33:37]
  wire [2:0] _T_642; // @[Lookup.scala 33:37]
  wire [2:0] _T_643; // @[Lookup.scala 33:37]
  wire [2:0] _T_644; // @[Lookup.scala 33:37]
  wire [2:0] _T_645; // @[Lookup.scala 33:37]
  wire [2:0] _T_646; // @[Lookup.scala 33:37]
  wire [2:0] _T_647; // @[Lookup.scala 33:37]
  wire [2:0] _T_648; // @[Lookup.scala 33:37]
  wire [2:0] _T_649; // @[Lookup.scala 33:37]
  wire [2:0] _T_650; // @[Lookup.scala 33:37]
  wire [2:0] _T_651; // @[Lookup.scala 33:37]
  wire [2:0] _T_652; // @[Lookup.scala 33:37]
  wire [2:0] _T_653; // @[Lookup.scala 33:37]
  wire [2:0] _T_654; // @[Lookup.scala 33:37]
  wire [2:0] _T_655; // @[Lookup.scala 33:37]
  wire [2:0] _T_656; // @[Lookup.scala 33:37]
  wire [2:0] _T_657; // @[Lookup.scala 33:37]
  wire [2:0] _T_658; // @[Lookup.scala 33:37]
  wire [2:0] _T_659; // @[Lookup.scala 33:37]
  wire [2:0] _T_660; // @[Lookup.scala 33:37]
  wire [2:0] _T_661; // @[Lookup.scala 33:37]
  wire [2:0] _T_662; // @[Lookup.scala 33:37]
  wire [2:0] _T_663; // @[Lookup.scala 33:37]
  wire [2:0] _T_664; // @[Lookup.scala 33:37]
  wire [2:0] _T_665; // @[Lookup.scala 33:37]
  wire [2:0] _T_666; // @[Lookup.scala 33:37]
  wire [2:0] _T_667; // @[Lookup.scala 33:37]
  wire [2:0] _T_668; // @[Lookup.scala 33:37]
  wire [2:0] _T_669; // @[Lookup.scala 33:37]
  wire [2:0] _T_670; // @[Lookup.scala 33:37]
  wire [2:0] _T_671; // @[Lookup.scala 33:37]
  wire [2:0] _T_672; // @[Lookup.scala 33:37]
  wire [2:0] _T_673; // @[Lookup.scala 33:37]
  wire  _T_674; // @[Lookup.scala 33:37]
  wire  _T_675; // @[Lookup.scala 33:37]
  wire  _T_676; // @[Lookup.scala 33:37]
  wire  _T_677; // @[Lookup.scala 33:37]
  wire  _T_678; // @[Lookup.scala 33:37]
  wire  _T_679; // @[Lookup.scala 33:37]
  wire  _T_680; // @[Lookup.scala 33:37]
  wire  _T_681; // @[Lookup.scala 33:37]
  wire  _T_682; // @[Lookup.scala 33:37]
  wire  _T_683; // @[Lookup.scala 33:37]
  wire  _T_684; // @[Lookup.scala 33:37]
  wire  _T_685; // @[Lookup.scala 33:37]
  wire  _T_686; // @[Lookup.scala 33:37]
  wire  _T_687; // @[Lookup.scala 33:37]
  wire  _T_688; // @[Lookup.scala 33:37]
  wire  _T_689; // @[Lookup.scala 33:37]
  wire  _T_690; // @[Lookup.scala 33:37]
  wire  _T_691; // @[Lookup.scala 33:37]
  wire  _T_692; // @[Lookup.scala 33:37]
  wire  _T_693; // @[Lookup.scala 33:37]
  wire  _T_694; // @[Lookup.scala 33:37]
  wire  _T_695; // @[Lookup.scala 33:37]
  wire  _T_696; // @[Lookup.scala 33:37]
  wire  _T_697; // @[Lookup.scala 33:37]
  wire  _T_698; // @[Lookup.scala 33:37]
  wire  _T_699; // @[Lookup.scala 33:37]
  wire  _T_700; // @[Lookup.scala 33:37]
  wire  _T_701; // @[Lookup.scala 33:37]
  wire  _T_702; // @[Lookup.scala 33:37]
  wire  _T_703; // @[Lookup.scala 33:37]
  wire  _T_704; // @[Lookup.scala 33:37]
  wire  _T_705; // @[Lookup.scala 33:37]
  wire  _T_706; // @[Lookup.scala 33:37]
  wire  _T_707; // @[Lookup.scala 33:37]
  wire  _T_708; // @[Lookup.scala 33:37]
  wire  _T_709; // @[Lookup.scala 33:37]
  wire  _T_710; // @[Lookup.scala 33:37]
  wire  _T_711; // @[Lookup.scala 33:37]
  wire  _T_712; // @[Lookup.scala 33:37]
  wire  _T_713; // @[Lookup.scala 33:37]
  wire  _T_714; // @[Lookup.scala 33:37]
  wire  _T_715; // @[Lookup.scala 33:37]
  wire  _T_716; // @[Lookup.scala 33:37]
  wire  _T_717; // @[Lookup.scala 33:37]
  wire  _T_718; // @[Lookup.scala 33:37]
  wire  _T_719; // @[Lookup.scala 33:37]
  wire  _T_720; // @[Lookup.scala 33:37]
  wire  _T_721; // @[Lookup.scala 33:37]
  assign _T = io_inst & 32'h7f; // @[Lookup.scala 31:38]
  assign _T_1 = 32'h37 == _T; // @[Lookup.scala 31:38]
  assign _T_3 = 32'h17 == _T; // @[Lookup.scala 31:38]
  assign _T_5 = 32'h6f == _T; // @[Lookup.scala 31:38]
  assign _T_6 = io_inst & 32'h707f; // @[Lookup.scala 31:38]
  assign _T_7 = 32'h67 == _T_6; // @[Lookup.scala 31:38]
  assign _T_9 = 32'h63 == _T_6; // @[Lookup.scala 31:38]
  assign _T_11 = 32'h1063 == _T_6; // @[Lookup.scala 31:38]
  assign _T_13 = 32'h4063 == _T_6; // @[Lookup.scala 31:38]
  assign _T_15 = 32'h5063 == _T_6; // @[Lookup.scala 31:38]
  assign _T_17 = 32'h6063 == _T_6; // @[Lookup.scala 31:38]
  assign _T_19 = 32'h7063 == _T_6; // @[Lookup.scala 31:38]
  assign _T_21 = 32'h3 == _T_6; // @[Lookup.scala 31:38]
  assign _T_23 = 32'h1003 == _T_6; // @[Lookup.scala 31:38]
  assign _T_25 = 32'h2003 == _T_6; // @[Lookup.scala 31:38]
  assign _T_27 = 32'h4003 == _T_6; // @[Lookup.scala 31:38]
  assign _T_29 = 32'h5003 == _T_6; // @[Lookup.scala 31:38]
  assign _T_31 = 32'h23 == _T_6; // @[Lookup.scala 31:38]
  assign _T_33 = 32'h1023 == _T_6; // @[Lookup.scala 31:38]
  assign _T_35 = 32'h2023 == _T_6; // @[Lookup.scala 31:38]
  assign _T_37 = 32'h13 == _T_6; // @[Lookup.scala 31:38]
  assign _T_39 = 32'h2013 == _T_6; // @[Lookup.scala 31:38]
  assign _T_41 = 32'h3013 == _T_6; // @[Lookup.scala 31:38]
  assign _T_43 = 32'h4013 == _T_6; // @[Lookup.scala 31:38]
  assign _T_45 = 32'h6013 == _T_6; // @[Lookup.scala 31:38]
  assign _T_47 = 32'h7013 == _T_6; // @[Lookup.scala 31:38]
  assign _T_48 = io_inst & 32'hfe00707f; // @[Lookup.scala 31:38]
  assign _T_49 = 32'h1013 == _T_48; // @[Lookup.scala 31:38]
  assign _T_51 = 32'h5013 == _T_48; // @[Lookup.scala 31:38]
  assign _T_53 = 32'h40005013 == _T_48; // @[Lookup.scala 31:38]
  assign _T_55 = 32'h33 == _T_48; // @[Lookup.scala 31:38]
  assign _T_57 = 32'h40000033 == _T_48; // @[Lookup.scala 31:38]
  assign _T_59 = 32'h1033 == _T_48; // @[Lookup.scala 31:38]
  assign _T_61 = 32'h2033 == _T_48; // @[Lookup.scala 31:38]
  assign _T_63 = 32'h3033 == _T_48; // @[Lookup.scala 31:38]
  assign _T_65 = 32'h4033 == _T_48; // @[Lookup.scala 31:38]
  assign _T_67 = 32'h5033 == _T_48; // @[Lookup.scala 31:38]
  assign _T_69 = 32'h40005033 == _T_48; // @[Lookup.scala 31:38]
  assign _T_71 = 32'h6033 == _T_48; // @[Lookup.scala 31:38]
  assign _T_73 = 32'h7033 == _T_48; // @[Lookup.scala 31:38]
  assign _T_74 = io_inst & 32'hf00fffff; // @[Lookup.scala 31:38]
  assign _T_75 = 32'hf == _T_74; // @[Lookup.scala 31:38]
  assign _T_77 = 32'h100f == io_inst; // @[Lookup.scala 31:38]
  assign _T_79 = 32'h1073 == _T_6; // @[Lookup.scala 31:38]
  assign _T_81 = 32'h2073 == _T_6; // @[Lookup.scala 31:38]
  assign _T_83 = 32'h3073 == _T_6; // @[Lookup.scala 31:38]
  assign _T_85 = 32'h5073 == _T_6; // @[Lookup.scala 31:38]
  assign _T_87 = 32'h6073 == _T_6; // @[Lookup.scala 31:38]
  assign _T_89 = 32'h7073 == _T_6; // @[Lookup.scala 31:38]
  assign _T_91 = 32'h73 == io_inst; // @[Lookup.scala 31:38]
  assign _T_93 = 32'h100073 == io_inst; // @[Lookup.scala 31:38]
  assign _T_95 = 32'h10000073 == io_inst; // @[Lookup.scala 31:38]
  assign _T_97 = 32'h10200073 == io_inst; // @[Lookup.scala 31:38]
  assign _T_99 = _T_95 ? 2'h3 : 2'h0; // @[Lookup.scala 33:37]
  assign _T_100 = _T_93 ? 2'h0 : _T_99; // @[Lookup.scala 33:37]
  assign _T_101 = _T_91 ? 2'h0 : _T_100; // @[Lookup.scala 33:37]
  assign _T_102 = _T_89 ? 2'h2 : _T_101; // @[Lookup.scala 33:37]
  assign _T_103 = _T_87 ? 2'h2 : _T_102; // @[Lookup.scala 33:37]
  assign _T_104 = _T_85 ? 2'h2 : _T_103; // @[Lookup.scala 33:37]
  assign _T_105 = _T_83 ? 2'h2 : _T_104; // @[Lookup.scala 33:37]
  assign _T_106 = _T_81 ? 2'h2 : _T_105; // @[Lookup.scala 33:37]
  assign _T_107 = _T_79 ? 2'h2 : _T_106; // @[Lookup.scala 33:37]
  assign _T_108 = _T_77 ? 2'h2 : _T_107; // @[Lookup.scala 33:37]
  assign _T_109 = _T_75 ? 2'h0 : _T_108; // @[Lookup.scala 33:37]
  assign _T_110 = _T_73 ? 2'h0 : _T_109; // @[Lookup.scala 33:37]
  assign _T_111 = _T_71 ? 2'h0 : _T_110; // @[Lookup.scala 33:37]
  assign _T_112 = _T_69 ? 2'h0 : _T_111; // @[Lookup.scala 33:37]
  assign _T_113 = _T_67 ? 2'h0 : _T_112; // @[Lookup.scala 33:37]
  assign _T_114 = _T_65 ? 2'h0 : _T_113; // @[Lookup.scala 33:37]
  assign _T_115 = _T_63 ? 2'h0 : _T_114; // @[Lookup.scala 33:37]
  assign _T_116 = _T_61 ? 2'h0 : _T_115; // @[Lookup.scala 33:37]
  assign _T_117 = _T_59 ? 2'h0 : _T_116; // @[Lookup.scala 33:37]
  assign _T_118 = _T_57 ? 2'h0 : _T_117; // @[Lookup.scala 33:37]
  assign _T_119 = _T_55 ? 2'h0 : _T_118; // @[Lookup.scala 33:37]
  assign _T_120 = _T_53 ? 2'h0 : _T_119; // @[Lookup.scala 33:37]
  assign _T_121 = _T_51 ? 2'h0 : _T_120; // @[Lookup.scala 33:37]
  assign _T_122 = _T_49 ? 2'h0 : _T_121; // @[Lookup.scala 33:37]
  assign _T_123 = _T_47 ? 2'h0 : _T_122; // @[Lookup.scala 33:37]
  assign _T_124 = _T_45 ? 2'h0 : _T_123; // @[Lookup.scala 33:37]
  assign _T_125 = _T_43 ? 2'h0 : _T_124; // @[Lookup.scala 33:37]
  assign _T_126 = _T_41 ? 2'h0 : _T_125; // @[Lookup.scala 33:37]
  assign _T_127 = _T_39 ? 2'h0 : _T_126; // @[Lookup.scala 33:37]
  assign _T_128 = _T_37 ? 2'h0 : _T_127; // @[Lookup.scala 33:37]
  assign _T_129 = _T_35 ? 2'h0 : _T_128; // @[Lookup.scala 33:37]
  assign _T_130 = _T_33 ? 2'h0 : _T_129; // @[Lookup.scala 33:37]
  assign _T_131 = _T_31 ? 2'h0 : _T_130; // @[Lookup.scala 33:37]
  assign _T_132 = _T_29 ? 2'h2 : _T_131; // @[Lookup.scala 33:37]
  assign _T_133 = _T_27 ? 2'h2 : _T_132; // @[Lookup.scala 33:37]
  assign _T_134 = _T_25 ? 2'h2 : _T_133; // @[Lookup.scala 33:37]
  assign _T_135 = _T_23 ? 2'h2 : _T_134; // @[Lookup.scala 33:37]
  assign _T_136 = _T_21 ? 2'h2 : _T_135; // @[Lookup.scala 33:37]
  assign _T_137 = _T_19 ? 2'h0 : _T_136; // @[Lookup.scala 33:37]
  assign _T_138 = _T_17 ? 2'h0 : _T_137; // @[Lookup.scala 33:37]
  assign _T_139 = _T_15 ? 2'h0 : _T_138; // @[Lookup.scala 33:37]
  assign _T_140 = _T_13 ? 2'h0 : _T_139; // @[Lookup.scala 33:37]
  assign _T_141 = _T_11 ? 2'h0 : _T_140; // @[Lookup.scala 33:37]
  assign _T_142 = _T_9 ? 2'h0 : _T_141; // @[Lookup.scala 33:37]
  assign _T_143 = _T_7 ? 2'h1 : _T_142; // @[Lookup.scala 33:37]
  assign _T_144 = _T_5 ? 2'h1 : _T_143; // @[Lookup.scala 33:37]
  assign _T_145 = _T_3 ? 2'h0 : _T_144; // @[Lookup.scala 33:37]
  assign _T_154 = _T_81 | _T_83; // @[Lookup.scala 33:37]
  assign _T_155 = _T_79 | _T_154; // @[Lookup.scala 33:37]
  assign _T_156 = _T_77 ? 1'h0 : _T_155; // @[Lookup.scala 33:37]
  assign _T_157 = _T_75 ? 1'h0 : _T_156; // @[Lookup.scala 33:37]
  assign _T_158 = _T_73 | _T_157; // @[Lookup.scala 33:37]
  assign _T_159 = _T_71 | _T_158; // @[Lookup.scala 33:37]
  assign _T_160 = _T_69 | _T_159; // @[Lookup.scala 33:37]
  assign _T_161 = _T_67 | _T_160; // @[Lookup.scala 33:37]
  assign _T_162 = _T_65 | _T_161; // @[Lookup.scala 33:37]
  assign _T_163 = _T_63 | _T_162; // @[Lookup.scala 33:37]
  assign _T_164 = _T_61 | _T_163; // @[Lookup.scala 33:37]
  assign _T_165 = _T_59 | _T_164; // @[Lookup.scala 33:37]
  assign _T_166 = _T_57 | _T_165; // @[Lookup.scala 33:37]
  assign _T_167 = _T_55 | _T_166; // @[Lookup.scala 33:37]
  assign _T_168 = _T_53 | _T_167; // @[Lookup.scala 33:37]
  assign _T_169 = _T_51 | _T_168; // @[Lookup.scala 33:37]
  assign _T_170 = _T_49 | _T_169; // @[Lookup.scala 33:37]
  assign _T_171 = _T_47 | _T_170; // @[Lookup.scala 33:37]
  assign _T_172 = _T_45 | _T_171; // @[Lookup.scala 33:37]
  assign _T_173 = _T_43 | _T_172; // @[Lookup.scala 33:37]
  assign _T_174 = _T_41 | _T_173; // @[Lookup.scala 33:37]
  assign _T_175 = _T_39 | _T_174; // @[Lookup.scala 33:37]
  assign _T_176 = _T_37 | _T_175; // @[Lookup.scala 33:37]
  assign _T_177 = _T_35 | _T_176; // @[Lookup.scala 33:37]
  assign _T_178 = _T_33 | _T_177; // @[Lookup.scala 33:37]
  assign _T_179 = _T_31 | _T_178; // @[Lookup.scala 33:37]
  assign _T_180 = _T_29 | _T_179; // @[Lookup.scala 33:37]
  assign _T_181 = _T_27 | _T_180; // @[Lookup.scala 33:37]
  assign _T_182 = _T_25 | _T_181; // @[Lookup.scala 33:37]
  assign _T_183 = _T_23 | _T_182; // @[Lookup.scala 33:37]
  assign _T_184 = _T_21 | _T_183; // @[Lookup.scala 33:37]
  assign _T_185 = _T_19 ? 1'h0 : _T_184; // @[Lookup.scala 33:37]
  assign _T_186 = _T_17 ? 1'h0 : _T_185; // @[Lookup.scala 33:37]
  assign _T_187 = _T_15 ? 1'h0 : _T_186; // @[Lookup.scala 33:37]
  assign _T_188 = _T_13 ? 1'h0 : _T_187; // @[Lookup.scala 33:37]
  assign _T_189 = _T_11 ? 1'h0 : _T_188; // @[Lookup.scala 33:37]
  assign _T_190 = _T_9 ? 1'h0 : _T_189; // @[Lookup.scala 33:37]
  assign _T_191 = _T_7 | _T_190; // @[Lookup.scala 33:37]
  assign _T_192 = _T_5 ? 1'h0 : _T_191; // @[Lookup.scala 33:37]
  assign _T_193 = _T_3 ? 1'h0 : _T_192; // @[Lookup.scala 33:37]
  assign _T_207 = _T_71 | _T_73; // @[Lookup.scala 33:37]
  assign _T_208 = _T_69 | _T_207; // @[Lookup.scala 33:37]
  assign _T_209 = _T_67 | _T_208; // @[Lookup.scala 33:37]
  assign _T_210 = _T_65 | _T_209; // @[Lookup.scala 33:37]
  assign _T_211 = _T_63 | _T_210; // @[Lookup.scala 33:37]
  assign _T_212 = _T_61 | _T_211; // @[Lookup.scala 33:37]
  assign _T_213 = _T_59 | _T_212; // @[Lookup.scala 33:37]
  assign _T_214 = _T_57 | _T_213; // @[Lookup.scala 33:37]
  assign _T_215 = _T_55 | _T_214; // @[Lookup.scala 33:37]
  assign _T_216 = _T_53 ? 1'h0 : _T_215; // @[Lookup.scala 33:37]
  assign _T_217 = _T_51 ? 1'h0 : _T_216; // @[Lookup.scala 33:37]
  assign _T_218 = _T_49 ? 1'h0 : _T_217; // @[Lookup.scala 33:37]
  assign _T_219 = _T_47 ? 1'h0 : _T_218; // @[Lookup.scala 33:37]
  assign _T_220 = _T_45 ? 1'h0 : _T_219; // @[Lookup.scala 33:37]
  assign _T_221 = _T_43 ? 1'h0 : _T_220; // @[Lookup.scala 33:37]
  assign _T_222 = _T_41 ? 1'h0 : _T_221; // @[Lookup.scala 33:37]
  assign _T_223 = _T_39 ? 1'h0 : _T_222; // @[Lookup.scala 33:37]
  assign _T_224 = _T_37 ? 1'h0 : _T_223; // @[Lookup.scala 33:37]
  assign _T_225 = _T_35 ? 1'h0 : _T_224; // @[Lookup.scala 33:37]
  assign _T_226 = _T_33 ? 1'h0 : _T_225; // @[Lookup.scala 33:37]
  assign _T_227 = _T_31 ? 1'h0 : _T_226; // @[Lookup.scala 33:37]
  assign _T_228 = _T_29 ? 1'h0 : _T_227; // @[Lookup.scala 33:37]
  assign _T_229 = _T_27 ? 1'h0 : _T_228; // @[Lookup.scala 33:37]
  assign _T_230 = _T_25 ? 1'h0 : _T_229; // @[Lookup.scala 33:37]
  assign _T_231 = _T_23 ? 1'h0 : _T_230; // @[Lookup.scala 33:37]
  assign _T_232 = _T_21 ? 1'h0 : _T_231; // @[Lookup.scala 33:37]
  assign _T_233 = _T_19 ? 1'h0 : _T_232; // @[Lookup.scala 33:37]
  assign _T_234 = _T_17 ? 1'h0 : _T_233; // @[Lookup.scala 33:37]
  assign _T_235 = _T_15 ? 1'h0 : _T_234; // @[Lookup.scala 33:37]
  assign _T_236 = _T_13 ? 1'h0 : _T_235; // @[Lookup.scala 33:37]
  assign _T_237 = _T_11 ? 1'h0 : _T_236; // @[Lookup.scala 33:37]
  assign _T_238 = _T_9 ? 1'h0 : _T_237; // @[Lookup.scala 33:37]
  assign _T_239 = _T_7 ? 1'h0 : _T_238; // @[Lookup.scala 33:37]
  assign _T_240 = _T_5 ? 1'h0 : _T_239; // @[Lookup.scala 33:37]
  assign _T_241 = _T_3 ? 1'h0 : _T_240; // @[Lookup.scala 33:37]
  assign _T_246 = _T_89 ? 3'h6 : 3'h0; // @[Lookup.scala 33:37]
  assign _T_247 = _T_87 ? 3'h6 : _T_246; // @[Lookup.scala 33:37]
  assign _T_248 = _T_85 ? 3'h6 : _T_247; // @[Lookup.scala 33:37]
  assign _T_249 = _T_83 ? 3'h0 : _T_248; // @[Lookup.scala 33:37]
  assign _T_250 = _T_81 ? 3'h0 : _T_249; // @[Lookup.scala 33:37]
  assign _T_251 = _T_79 ? 3'h0 : _T_250; // @[Lookup.scala 33:37]
  assign _T_252 = _T_77 ? 3'h0 : _T_251; // @[Lookup.scala 33:37]
  assign _T_253 = _T_75 ? 3'h0 : _T_252; // @[Lookup.scala 33:37]
  assign _T_254 = _T_73 ? 3'h0 : _T_253; // @[Lookup.scala 33:37]
  assign _T_255 = _T_71 ? 3'h0 : _T_254; // @[Lookup.scala 33:37]
  assign _T_256 = _T_69 ? 3'h0 : _T_255; // @[Lookup.scala 33:37]
  assign _T_257 = _T_67 ? 3'h0 : _T_256; // @[Lookup.scala 33:37]
  assign _T_258 = _T_65 ? 3'h0 : _T_257; // @[Lookup.scala 33:37]
  assign _T_259 = _T_63 ? 3'h0 : _T_258; // @[Lookup.scala 33:37]
  assign _T_260 = _T_61 ? 3'h0 : _T_259; // @[Lookup.scala 33:37]
  assign _T_261 = _T_59 ? 3'h0 : _T_260; // @[Lookup.scala 33:37]
  assign _T_262 = _T_57 ? 3'h0 : _T_261; // @[Lookup.scala 33:37]
  assign _T_263 = _T_55 ? 3'h0 : _T_262; // @[Lookup.scala 33:37]
  assign _T_264 = _T_53 ? 3'h1 : _T_263; // @[Lookup.scala 33:37]
  assign _T_265 = _T_51 ? 3'h1 : _T_264; // @[Lookup.scala 33:37]
  assign _T_266 = _T_49 ? 3'h1 : _T_265; // @[Lookup.scala 33:37]
  assign _T_267 = _T_47 ? 3'h1 : _T_266; // @[Lookup.scala 33:37]
  assign _T_268 = _T_45 ? 3'h1 : _T_267; // @[Lookup.scala 33:37]
  assign _T_269 = _T_43 ? 3'h1 : _T_268; // @[Lookup.scala 33:37]
  assign _T_270 = _T_41 ? 3'h1 : _T_269; // @[Lookup.scala 33:37]
  assign _T_271 = _T_39 ? 3'h1 : _T_270; // @[Lookup.scala 33:37]
  assign _T_272 = _T_37 ? 3'h1 : _T_271; // @[Lookup.scala 33:37]
  assign _T_273 = _T_35 ? 3'h2 : _T_272; // @[Lookup.scala 33:37]
  assign _T_274 = _T_33 ? 3'h2 : _T_273; // @[Lookup.scala 33:37]
  assign _T_275 = _T_31 ? 3'h2 : _T_274; // @[Lookup.scala 33:37]
  assign _T_276 = _T_29 ? 3'h1 : _T_275; // @[Lookup.scala 33:37]
  assign _T_277 = _T_27 ? 3'h1 : _T_276; // @[Lookup.scala 33:37]
  assign _T_278 = _T_25 ? 3'h1 : _T_277; // @[Lookup.scala 33:37]
  assign _T_279 = _T_23 ? 3'h1 : _T_278; // @[Lookup.scala 33:37]
  assign _T_280 = _T_21 ? 3'h1 : _T_279; // @[Lookup.scala 33:37]
  assign _T_281 = _T_19 ? 3'h5 : _T_280; // @[Lookup.scala 33:37]
  assign _T_282 = _T_17 ? 3'h5 : _T_281; // @[Lookup.scala 33:37]
  assign _T_283 = _T_15 ? 3'h5 : _T_282; // @[Lookup.scala 33:37]
  assign _T_284 = _T_13 ? 3'h5 : _T_283; // @[Lookup.scala 33:37]
  assign _T_285 = _T_11 ? 3'h5 : _T_284; // @[Lookup.scala 33:37]
  assign _T_286 = _T_9 ? 3'h5 : _T_285; // @[Lookup.scala 33:37]
  assign _T_287 = _T_7 ? 3'h1 : _T_286; // @[Lookup.scala 33:37]
  assign _T_288 = _T_5 ? 3'h4 : _T_287; // @[Lookup.scala 33:37]
  assign _T_289 = _T_3 ? 3'h3 : _T_288; // @[Lookup.scala 33:37]
  assign _T_297 = _T_83 ? 4'ha : 4'hf; // @[Lookup.scala 33:37]
  assign _T_298 = _T_81 ? 4'ha : _T_297; // @[Lookup.scala 33:37]
  assign _T_299 = _T_79 ? 4'ha : _T_298; // @[Lookup.scala 33:37]
  assign _T_300 = _T_77 ? 4'hf : _T_299; // @[Lookup.scala 33:37]
  assign _T_301 = _T_75 ? 4'hf : _T_300; // @[Lookup.scala 33:37]
  assign _T_302 = _T_73 ? 4'h2 : _T_301; // @[Lookup.scala 33:37]
  assign _T_303 = _T_71 ? 4'h3 : _T_302; // @[Lookup.scala 33:37]
  assign _T_304 = _T_69 ? 4'h9 : _T_303; // @[Lookup.scala 33:37]
  assign _T_305 = _T_67 ? 4'h8 : _T_304; // @[Lookup.scala 33:37]
  assign _T_306 = _T_65 ? 4'h4 : _T_305; // @[Lookup.scala 33:37]
  assign _T_307 = _T_63 ? 4'h7 : _T_306; // @[Lookup.scala 33:37]
  assign _T_308 = _T_61 ? 4'h5 : _T_307; // @[Lookup.scala 33:37]
  assign _T_309 = _T_59 ? 4'h6 : _T_308; // @[Lookup.scala 33:37]
  assign _T_310 = _T_57 ? 4'h1 : _T_309; // @[Lookup.scala 33:37]
  assign _T_311 = _T_55 ? 4'h0 : _T_310; // @[Lookup.scala 33:37]
  assign _T_312 = _T_53 ? 4'h9 : _T_311; // @[Lookup.scala 33:37]
  assign _T_313 = _T_51 ? 4'h8 : _T_312; // @[Lookup.scala 33:37]
  assign _T_314 = _T_49 ? 4'h6 : _T_313; // @[Lookup.scala 33:37]
  assign _T_315 = _T_47 ? 4'h2 : _T_314; // @[Lookup.scala 33:37]
  assign _T_316 = _T_45 ? 4'h3 : _T_315; // @[Lookup.scala 33:37]
  assign _T_317 = _T_43 ? 4'h4 : _T_316; // @[Lookup.scala 33:37]
  assign _T_318 = _T_41 ? 4'h7 : _T_317; // @[Lookup.scala 33:37]
  assign _T_319 = _T_39 ? 4'h5 : _T_318; // @[Lookup.scala 33:37]
  assign _T_320 = _T_37 ? 4'h0 : _T_319; // @[Lookup.scala 33:37]
  assign _T_321 = _T_35 ? 4'h0 : _T_320; // @[Lookup.scala 33:37]
  assign _T_322 = _T_33 ? 4'h0 : _T_321; // @[Lookup.scala 33:37]
  assign _T_323 = _T_31 ? 4'h0 : _T_322; // @[Lookup.scala 33:37]
  assign _T_324 = _T_29 ? 4'h0 : _T_323; // @[Lookup.scala 33:37]
  assign _T_325 = _T_27 ? 4'h0 : _T_324; // @[Lookup.scala 33:37]
  assign _T_326 = _T_25 ? 4'h0 : _T_325; // @[Lookup.scala 33:37]
  assign _T_327 = _T_23 ? 4'h0 : _T_326; // @[Lookup.scala 33:37]
  assign _T_328 = _T_21 ? 4'h0 : _T_327; // @[Lookup.scala 33:37]
  assign _T_329 = _T_19 ? 4'h0 : _T_328; // @[Lookup.scala 33:37]
  assign _T_330 = _T_17 ? 4'h0 : _T_329; // @[Lookup.scala 33:37]
  assign _T_331 = _T_15 ? 4'h0 : _T_330; // @[Lookup.scala 33:37]
  assign _T_332 = _T_13 ? 4'h0 : _T_331; // @[Lookup.scala 33:37]
  assign _T_333 = _T_11 ? 4'h0 : _T_332; // @[Lookup.scala 33:37]
  assign _T_334 = _T_9 ? 4'h0 : _T_333; // @[Lookup.scala 33:37]
  assign _T_335 = _T_7 ? 4'h0 : _T_334; // @[Lookup.scala 33:37]
  assign _T_336 = _T_5 ? 4'h0 : _T_335; // @[Lookup.scala 33:37]
  assign _T_337 = _T_3 ? 4'h0 : _T_336; // @[Lookup.scala 33:37]
  assign _T_377 = _T_19 ? 3'h4 : 3'h0; // @[Lookup.scala 33:37]
  assign _T_378 = _T_17 ? 3'h1 : _T_377; // @[Lookup.scala 33:37]
  assign _T_379 = _T_15 ? 3'h5 : _T_378; // @[Lookup.scala 33:37]
  assign _T_380 = _T_13 ? 3'h2 : _T_379; // @[Lookup.scala 33:37]
  assign _T_381 = _T_11 ? 3'h6 : _T_380; // @[Lookup.scala 33:37]
  assign _T_382 = _T_9 ? 3'h3 : _T_381; // @[Lookup.scala 33:37]
  assign _T_383 = _T_7 ? 3'h0 : _T_382; // @[Lookup.scala 33:37]
  assign _T_384 = _T_5 ? 3'h0 : _T_383; // @[Lookup.scala 33:37]
  assign _T_385 = _T_3 ? 3'h0 : _T_384; // @[Lookup.scala 33:37]
  assign _T_388 = _T_93 ? 1'h0 : _T_95; // @[Lookup.scala 33:37]
  assign _T_389 = _T_91 ? 1'h0 : _T_388; // @[Lookup.scala 33:37]
  assign _T_390 = _T_89 | _T_389; // @[Lookup.scala 33:37]
  assign _T_391 = _T_87 | _T_390; // @[Lookup.scala 33:37]
  assign _T_392 = _T_85 | _T_391; // @[Lookup.scala 33:37]
  assign _T_393 = _T_83 | _T_392; // @[Lookup.scala 33:37]
  assign _T_394 = _T_81 | _T_393; // @[Lookup.scala 33:37]
  assign _T_395 = _T_79 | _T_394; // @[Lookup.scala 33:37]
  assign _T_396 = _T_77 | _T_395; // @[Lookup.scala 33:37]
  assign _T_397 = _T_75 ? 1'h0 : _T_396; // @[Lookup.scala 33:37]
  assign _T_398 = _T_73 ? 1'h0 : _T_397; // @[Lookup.scala 33:37]
  assign _T_399 = _T_71 ? 1'h0 : _T_398; // @[Lookup.scala 33:37]
  assign _T_400 = _T_69 ? 1'h0 : _T_399; // @[Lookup.scala 33:37]
  assign _T_401 = _T_67 ? 1'h0 : _T_400; // @[Lookup.scala 33:37]
  assign _T_402 = _T_65 ? 1'h0 : _T_401; // @[Lookup.scala 33:37]
  assign _T_403 = _T_63 ? 1'h0 : _T_402; // @[Lookup.scala 33:37]
  assign _T_404 = _T_61 ? 1'h0 : _T_403; // @[Lookup.scala 33:37]
  assign _T_405 = _T_59 ? 1'h0 : _T_404; // @[Lookup.scala 33:37]
  assign _T_406 = _T_57 ? 1'h0 : _T_405; // @[Lookup.scala 33:37]
  assign _T_407 = _T_55 ? 1'h0 : _T_406; // @[Lookup.scala 33:37]
  assign _T_408 = _T_53 ? 1'h0 : _T_407; // @[Lookup.scala 33:37]
  assign _T_409 = _T_51 ? 1'h0 : _T_408; // @[Lookup.scala 33:37]
  assign _T_410 = _T_49 ? 1'h0 : _T_409; // @[Lookup.scala 33:37]
  assign _T_411 = _T_47 ? 1'h0 : _T_410; // @[Lookup.scala 33:37]
  assign _T_412 = _T_45 ? 1'h0 : _T_411; // @[Lookup.scala 33:37]
  assign _T_413 = _T_43 ? 1'h0 : _T_412; // @[Lookup.scala 33:37]
  assign _T_414 = _T_41 ? 1'h0 : _T_413; // @[Lookup.scala 33:37]
  assign _T_415 = _T_39 ? 1'h0 : _T_414; // @[Lookup.scala 33:37]
  assign _T_416 = _T_37 ? 1'h0 : _T_415; // @[Lookup.scala 33:37]
  assign _T_417 = _T_35 ? 1'h0 : _T_416; // @[Lookup.scala 33:37]
  assign _T_418 = _T_33 ? 1'h0 : _T_417; // @[Lookup.scala 33:37]
  assign _T_419 = _T_31 ? 1'h0 : _T_418; // @[Lookup.scala 33:37]
  assign _T_420 = _T_29 | _T_419; // @[Lookup.scala 33:37]
  assign _T_421 = _T_27 | _T_420; // @[Lookup.scala 33:37]
  assign _T_422 = _T_25 | _T_421; // @[Lookup.scala 33:37]
  assign _T_423 = _T_23 | _T_422; // @[Lookup.scala 33:37]
  assign _T_424 = _T_21 | _T_423; // @[Lookup.scala 33:37]
  assign _T_425 = _T_19 ? 1'h0 : _T_424; // @[Lookup.scala 33:37]
  assign _T_426 = _T_17 ? 1'h0 : _T_425; // @[Lookup.scala 33:37]
  assign _T_427 = _T_15 ? 1'h0 : _T_426; // @[Lookup.scala 33:37]
  assign _T_428 = _T_13 ? 1'h0 : _T_427; // @[Lookup.scala 33:37]
  assign _T_429 = _T_11 ? 1'h0 : _T_428; // @[Lookup.scala 33:37]
  assign _T_430 = _T_9 ? 1'h0 : _T_429; // @[Lookup.scala 33:37]
  assign _T_431 = _T_7 | _T_430; // @[Lookup.scala 33:37]
  assign _T_432 = _T_5 | _T_431; // @[Lookup.scala 33:37]
  assign _T_433 = _T_3 ? 1'h0 : _T_432; // @[Lookup.scala 33:37]
  assign _T_465 = _T_35 ? 2'h1 : 2'h0; // @[Lookup.scala 33:37]
  assign _T_466 = _T_33 ? 2'h2 : _T_465; // @[Lookup.scala 33:37]
  assign _T_467 = _T_31 ? 2'h3 : _T_466; // @[Lookup.scala 33:37]
  assign _T_468 = _T_29 ? 2'h0 : _T_467; // @[Lookup.scala 33:37]
  assign _T_469 = _T_27 ? 2'h0 : _T_468; // @[Lookup.scala 33:37]
  assign _T_470 = _T_25 ? 2'h0 : _T_469; // @[Lookup.scala 33:37]
  assign _T_471 = _T_23 ? 2'h0 : _T_470; // @[Lookup.scala 33:37]
  assign _T_472 = _T_21 ? 2'h0 : _T_471; // @[Lookup.scala 33:37]
  assign _T_473 = _T_19 ? 2'h0 : _T_472; // @[Lookup.scala 33:37]
  assign _T_474 = _T_17 ? 2'h0 : _T_473; // @[Lookup.scala 33:37]
  assign _T_475 = _T_15 ? 2'h0 : _T_474; // @[Lookup.scala 33:37]
  assign _T_476 = _T_13 ? 2'h0 : _T_475; // @[Lookup.scala 33:37]
  assign _T_477 = _T_11 ? 2'h0 : _T_476; // @[Lookup.scala 33:37]
  assign _T_478 = _T_9 ? 2'h0 : _T_477; // @[Lookup.scala 33:37]
  assign _T_479 = _T_7 ? 2'h0 : _T_478; // @[Lookup.scala 33:37]
  assign _T_480 = _T_5 ? 2'h0 : _T_479; // @[Lookup.scala 33:37]
  assign _T_481 = _T_3 ? 2'h0 : _T_480; // @[Lookup.scala 33:37]
  assign _T_516 = _T_29 ? 3'h4 : 3'h0; // @[Lookup.scala 33:37]
  assign _T_517 = _T_27 ? 3'h5 : _T_516; // @[Lookup.scala 33:37]
  assign _T_518 = _T_25 ? 3'h1 : _T_517; // @[Lookup.scala 33:37]
  assign _T_519 = _T_23 ? 3'h2 : _T_518; // @[Lookup.scala 33:37]
  assign _T_520 = _T_21 ? 3'h3 : _T_519; // @[Lookup.scala 33:37]
  assign _T_521 = _T_19 ? 3'h0 : _T_520; // @[Lookup.scala 33:37]
  assign _T_522 = _T_17 ? 3'h0 : _T_521; // @[Lookup.scala 33:37]
  assign _T_523 = _T_15 ? 3'h0 : _T_522; // @[Lookup.scala 33:37]
  assign _T_524 = _T_13 ? 3'h0 : _T_523; // @[Lookup.scala 33:37]
  assign _T_525 = _T_11 ? 3'h0 : _T_524; // @[Lookup.scala 33:37]
  assign _T_526 = _T_9 ? 3'h0 : _T_525; // @[Lookup.scala 33:37]
  assign _T_527 = _T_7 ? 3'h0 : _T_526; // @[Lookup.scala 33:37]
  assign _T_528 = _T_5 ? 3'h0 : _T_527; // @[Lookup.scala 33:37]
  assign _T_529 = _T_3 ? 3'h0 : _T_528; // @[Lookup.scala 33:37]
  assign _T_532 = _T_93 ? 2'h3 : _T_99; // @[Lookup.scala 33:37]
  assign _T_533 = _T_91 ? 2'h3 : _T_532; // @[Lookup.scala 33:37]
  assign _T_534 = _T_89 ? 2'h3 : _T_533; // @[Lookup.scala 33:37]
  assign _T_535 = _T_87 ? 2'h3 : _T_534; // @[Lookup.scala 33:37]
  assign _T_536 = _T_85 ? 2'h3 : _T_535; // @[Lookup.scala 33:37]
  assign _T_537 = _T_83 ? 2'h3 : _T_536; // @[Lookup.scala 33:37]
  assign _T_538 = _T_81 ? 2'h3 : _T_537; // @[Lookup.scala 33:37]
  assign _T_539 = _T_79 ? 2'h3 : _T_538; // @[Lookup.scala 33:37]
  assign _T_540 = _T_77 ? 2'h0 : _T_539; // @[Lookup.scala 33:37]
  assign _T_541 = _T_75 ? 2'h0 : _T_540; // @[Lookup.scala 33:37]
  assign _T_542 = _T_73 ? 2'h0 : _T_541; // @[Lookup.scala 33:37]
  assign _T_543 = _T_71 ? 2'h0 : _T_542; // @[Lookup.scala 33:37]
  assign _T_544 = _T_69 ? 2'h0 : _T_543; // @[Lookup.scala 33:37]
  assign _T_545 = _T_67 ? 2'h0 : _T_544; // @[Lookup.scala 33:37]
  assign _T_546 = _T_65 ? 2'h0 : _T_545; // @[Lookup.scala 33:37]
  assign _T_547 = _T_63 ? 2'h0 : _T_546; // @[Lookup.scala 33:37]
  assign _T_548 = _T_61 ? 2'h0 : _T_547; // @[Lookup.scala 33:37]
  assign _T_549 = _T_59 ? 2'h0 : _T_548; // @[Lookup.scala 33:37]
  assign _T_550 = _T_57 ? 2'h0 : _T_549; // @[Lookup.scala 33:37]
  assign _T_551 = _T_55 ? 2'h0 : _T_550; // @[Lookup.scala 33:37]
  assign _T_552 = _T_53 ? 2'h0 : _T_551; // @[Lookup.scala 33:37]
  assign _T_553 = _T_51 ? 2'h0 : _T_552; // @[Lookup.scala 33:37]
  assign _T_554 = _T_49 ? 2'h0 : _T_553; // @[Lookup.scala 33:37]
  assign _T_555 = _T_47 ? 2'h0 : _T_554; // @[Lookup.scala 33:37]
  assign _T_556 = _T_45 ? 2'h0 : _T_555; // @[Lookup.scala 33:37]
  assign _T_557 = _T_43 ? 2'h0 : _T_556; // @[Lookup.scala 33:37]
  assign _T_558 = _T_41 ? 2'h0 : _T_557; // @[Lookup.scala 33:37]
  assign _T_559 = _T_39 ? 2'h0 : _T_558; // @[Lookup.scala 33:37]
  assign _T_560 = _T_37 ? 2'h0 : _T_559; // @[Lookup.scala 33:37]
  assign _T_561 = _T_35 ? 2'h0 : _T_560; // @[Lookup.scala 33:37]
  assign _T_562 = _T_33 ? 2'h0 : _T_561; // @[Lookup.scala 33:37]
  assign _T_563 = _T_31 ? 2'h0 : _T_562; // @[Lookup.scala 33:37]
  assign _T_564 = _T_29 ? 2'h1 : _T_563; // @[Lookup.scala 33:37]
  assign _T_565 = _T_27 ? 2'h1 : _T_564; // @[Lookup.scala 33:37]
  assign _T_566 = _T_25 ? 2'h1 : _T_565; // @[Lookup.scala 33:37]
  assign _T_567 = _T_23 ? 2'h1 : _T_566; // @[Lookup.scala 33:37]
  assign _T_568 = _T_21 ? 2'h1 : _T_567; // @[Lookup.scala 33:37]
  assign _T_569 = _T_19 ? 2'h0 : _T_568; // @[Lookup.scala 33:37]
  assign _T_570 = _T_17 ? 2'h0 : _T_569; // @[Lookup.scala 33:37]
  assign _T_571 = _T_15 ? 2'h0 : _T_570; // @[Lookup.scala 33:37]
  assign _T_572 = _T_13 ? 2'h0 : _T_571; // @[Lookup.scala 33:37]
  assign _T_573 = _T_11 ? 2'h0 : _T_572; // @[Lookup.scala 33:37]
  assign _T_574 = _T_9 ? 2'h0 : _T_573; // @[Lookup.scala 33:37]
  assign _T_575 = _T_7 ? 2'h2 : _T_574; // @[Lookup.scala 33:37]
  assign _T_576 = _T_5 ? 2'h2 : _T_575; // @[Lookup.scala 33:37]
  assign _T_577 = _T_3 ? 2'h0 : _T_576; // @[Lookup.scala 33:37]
  assign _T_583 = _T_87 | _T_89; // @[Lookup.scala 33:37]
  assign _T_584 = _T_85 | _T_583; // @[Lookup.scala 33:37]
  assign _T_585 = _T_83 | _T_584; // @[Lookup.scala 33:37]
  assign _T_586 = _T_81 | _T_585; // @[Lookup.scala 33:37]
  assign _T_587 = _T_79 | _T_586; // @[Lookup.scala 33:37]
  assign _T_588 = _T_77 ? 1'h0 : _T_587; // @[Lookup.scala 33:37]
  assign _T_589 = _T_75 ? 1'h0 : _T_588; // @[Lookup.scala 33:37]
  assign _T_590 = _T_73 | _T_589; // @[Lookup.scala 33:37]
  assign _T_591 = _T_71 | _T_590; // @[Lookup.scala 33:37]
  assign _T_592 = _T_69 | _T_591; // @[Lookup.scala 33:37]
  assign _T_593 = _T_67 | _T_592; // @[Lookup.scala 33:37]
  assign _T_594 = _T_65 | _T_593; // @[Lookup.scala 33:37]
  assign _T_595 = _T_63 | _T_594; // @[Lookup.scala 33:37]
  assign _T_596 = _T_61 | _T_595; // @[Lookup.scala 33:37]
  assign _T_597 = _T_59 | _T_596; // @[Lookup.scala 33:37]
  assign _T_598 = _T_57 | _T_597; // @[Lookup.scala 33:37]
  assign _T_599 = _T_55 | _T_598; // @[Lookup.scala 33:37]
  assign _T_600 = _T_53 | _T_599; // @[Lookup.scala 33:37]
  assign _T_601 = _T_51 | _T_600; // @[Lookup.scala 33:37]
  assign _T_602 = _T_49 | _T_601; // @[Lookup.scala 33:37]
  assign _T_603 = _T_47 | _T_602; // @[Lookup.scala 33:37]
  assign _T_604 = _T_45 | _T_603; // @[Lookup.scala 33:37]
  assign _T_605 = _T_43 | _T_604; // @[Lookup.scala 33:37]
  assign _T_606 = _T_41 | _T_605; // @[Lookup.scala 33:37]
  assign _T_607 = _T_39 | _T_606; // @[Lookup.scala 33:37]
  assign _T_608 = _T_37 | _T_607; // @[Lookup.scala 33:37]
  assign _T_609 = _T_35 ? 1'h0 : _T_608; // @[Lookup.scala 33:37]
  assign _T_610 = _T_33 ? 1'h0 : _T_609; // @[Lookup.scala 33:37]
  assign _T_611 = _T_31 ? 1'h0 : _T_610; // @[Lookup.scala 33:37]
  assign _T_612 = _T_29 | _T_611; // @[Lookup.scala 33:37]
  assign _T_613 = _T_27 | _T_612; // @[Lookup.scala 33:37]
  assign _T_614 = _T_25 | _T_613; // @[Lookup.scala 33:37]
  assign _T_615 = _T_23 | _T_614; // @[Lookup.scala 33:37]
  assign _T_616 = _T_21 | _T_615; // @[Lookup.scala 33:37]
  assign _T_617 = _T_19 ? 1'h0 : _T_616; // @[Lookup.scala 33:37]
  assign _T_618 = _T_17 ? 1'h0 : _T_617; // @[Lookup.scala 33:37]
  assign _T_619 = _T_15 ? 1'h0 : _T_618; // @[Lookup.scala 33:37]
  assign _T_620 = _T_13 ? 1'h0 : _T_619; // @[Lookup.scala 33:37]
  assign _T_621 = _T_11 ? 1'h0 : _T_620; // @[Lookup.scala 33:37]
  assign _T_622 = _T_9 ? 1'h0 : _T_621; // @[Lookup.scala 33:37]
  assign _T_623 = _T_7 | _T_622; // @[Lookup.scala 33:37]
  assign _T_624 = _T_5 | _T_623; // @[Lookup.scala 33:37]
  assign _T_625 = _T_3 | _T_624; // @[Lookup.scala 33:37]
  assign _T_627 = _T_95 ? 3'h4 : 3'h0; // @[Lookup.scala 33:37]
  assign _T_628 = _T_93 ? 3'h4 : _T_627; // @[Lookup.scala 33:37]
  assign _T_629 = _T_91 ? 3'h4 : _T_628; // @[Lookup.scala 33:37]
  assign _T_630 = _T_89 ? 3'h3 : _T_629; // @[Lookup.scala 33:37]
  assign _T_631 = _T_87 ? 3'h2 : _T_630; // @[Lookup.scala 33:37]
  assign _T_632 = _T_85 ? 3'h1 : _T_631; // @[Lookup.scala 33:37]
  assign _T_633 = _T_83 ? 3'h3 : _T_632; // @[Lookup.scala 33:37]
  assign _T_634 = _T_81 ? 3'h2 : _T_633; // @[Lookup.scala 33:37]
  assign _T_635 = _T_79 ? 3'h1 : _T_634; // @[Lookup.scala 33:37]
  assign _T_636 = _T_77 ? 3'h0 : _T_635; // @[Lookup.scala 33:37]
  assign _T_637 = _T_75 ? 3'h0 : _T_636; // @[Lookup.scala 33:37]
  assign _T_638 = _T_73 ? 3'h0 : _T_637; // @[Lookup.scala 33:37]
  assign _T_639 = _T_71 ? 3'h0 : _T_638; // @[Lookup.scala 33:37]
  assign _T_640 = _T_69 ? 3'h0 : _T_639; // @[Lookup.scala 33:37]
  assign _T_641 = _T_67 ? 3'h0 : _T_640; // @[Lookup.scala 33:37]
  assign _T_642 = _T_65 ? 3'h0 : _T_641; // @[Lookup.scala 33:37]
  assign _T_643 = _T_63 ? 3'h0 : _T_642; // @[Lookup.scala 33:37]
  assign _T_644 = _T_61 ? 3'h0 : _T_643; // @[Lookup.scala 33:37]
  assign _T_645 = _T_59 ? 3'h0 : _T_644; // @[Lookup.scala 33:37]
  assign _T_646 = _T_57 ? 3'h0 : _T_645; // @[Lookup.scala 33:37]
  assign _T_647 = _T_55 ? 3'h0 : _T_646; // @[Lookup.scala 33:37]
  assign _T_648 = _T_53 ? 3'h0 : _T_647; // @[Lookup.scala 33:37]
  assign _T_649 = _T_51 ? 3'h0 : _T_648; // @[Lookup.scala 33:37]
  assign _T_650 = _T_49 ? 3'h0 : _T_649; // @[Lookup.scala 33:37]
  assign _T_651 = _T_47 ? 3'h0 : _T_650; // @[Lookup.scala 33:37]
  assign _T_652 = _T_45 ? 3'h0 : _T_651; // @[Lookup.scala 33:37]
  assign _T_653 = _T_43 ? 3'h0 : _T_652; // @[Lookup.scala 33:37]
  assign _T_654 = _T_41 ? 3'h0 : _T_653; // @[Lookup.scala 33:37]
  assign _T_655 = _T_39 ? 3'h0 : _T_654; // @[Lookup.scala 33:37]
  assign _T_656 = _T_37 ? 3'h0 : _T_655; // @[Lookup.scala 33:37]
  assign _T_657 = _T_35 ? 3'h0 : _T_656; // @[Lookup.scala 33:37]
  assign _T_658 = _T_33 ? 3'h0 : _T_657; // @[Lookup.scala 33:37]
  assign _T_659 = _T_31 ? 3'h0 : _T_658; // @[Lookup.scala 33:37]
  assign _T_660 = _T_29 ? 3'h0 : _T_659; // @[Lookup.scala 33:37]
  assign _T_661 = _T_27 ? 3'h0 : _T_660; // @[Lookup.scala 33:37]
  assign _T_662 = _T_25 ? 3'h0 : _T_661; // @[Lookup.scala 33:37]
  assign _T_663 = _T_23 ? 3'h0 : _T_662; // @[Lookup.scala 33:37]
  assign _T_664 = _T_21 ? 3'h0 : _T_663; // @[Lookup.scala 33:37]
  assign _T_665 = _T_19 ? 3'h0 : _T_664; // @[Lookup.scala 33:37]
  assign _T_666 = _T_17 ? 3'h0 : _T_665; // @[Lookup.scala 33:37]
  assign _T_667 = _T_15 ? 3'h0 : _T_666; // @[Lookup.scala 33:37]
  assign _T_668 = _T_13 ? 3'h0 : _T_667; // @[Lookup.scala 33:37]
  assign _T_669 = _T_11 ? 3'h0 : _T_668; // @[Lookup.scala 33:37]
  assign _T_670 = _T_9 ? 3'h0 : _T_669; // @[Lookup.scala 33:37]
  assign _T_671 = _T_7 ? 3'h0 : _T_670; // @[Lookup.scala 33:37]
  assign _T_672 = _T_5 ? 3'h0 : _T_671; // @[Lookup.scala 33:37]
  assign _T_673 = _T_3 ? 3'h0 : _T_672; // @[Lookup.scala 33:37]
  assign _T_674 = _T_97 ? 1'h0 : 1'h1; // @[Lookup.scala 33:37]
  assign _T_675 = _T_95 ? 1'h0 : _T_674; // @[Lookup.scala 33:37]
  assign _T_676 = _T_93 ? 1'h0 : _T_675; // @[Lookup.scala 33:37]
  assign _T_677 = _T_91 ? 1'h0 : _T_676; // @[Lookup.scala 33:37]
  assign _T_678 = _T_89 ? 1'h0 : _T_677; // @[Lookup.scala 33:37]
  assign _T_679 = _T_87 ? 1'h0 : _T_678; // @[Lookup.scala 33:37]
  assign _T_680 = _T_85 ? 1'h0 : _T_679; // @[Lookup.scala 33:37]
  assign _T_681 = _T_83 ? 1'h0 : _T_680; // @[Lookup.scala 33:37]
  assign _T_682 = _T_81 ? 1'h0 : _T_681; // @[Lookup.scala 33:37]
  assign _T_683 = _T_79 ? 1'h0 : _T_682; // @[Lookup.scala 33:37]
  assign _T_684 = _T_77 ? 1'h0 : _T_683; // @[Lookup.scala 33:37]
  assign _T_685 = _T_75 ? 1'h0 : _T_684; // @[Lookup.scala 33:37]
  assign _T_686 = _T_73 ? 1'h0 : _T_685; // @[Lookup.scala 33:37]
  assign _T_687 = _T_71 ? 1'h0 : _T_686; // @[Lookup.scala 33:37]
  assign _T_688 = _T_69 ? 1'h0 : _T_687; // @[Lookup.scala 33:37]
  assign _T_689 = _T_67 ? 1'h0 : _T_688; // @[Lookup.scala 33:37]
  assign _T_690 = _T_65 ? 1'h0 : _T_689; // @[Lookup.scala 33:37]
  assign _T_691 = _T_63 ? 1'h0 : _T_690; // @[Lookup.scala 33:37]
  assign _T_692 = _T_61 ? 1'h0 : _T_691; // @[Lookup.scala 33:37]
  assign _T_693 = _T_59 ? 1'h0 : _T_692; // @[Lookup.scala 33:37]
  assign _T_694 = _T_57 ? 1'h0 : _T_693; // @[Lookup.scala 33:37]
  assign _T_695 = _T_55 ? 1'h0 : _T_694; // @[Lookup.scala 33:37]
  assign _T_696 = _T_53 ? 1'h0 : _T_695; // @[Lookup.scala 33:37]
  assign _T_697 = _T_51 ? 1'h0 : _T_696; // @[Lookup.scala 33:37]
  assign _T_698 = _T_49 ? 1'h0 : _T_697; // @[Lookup.scala 33:37]
  assign _T_699 = _T_47 ? 1'h0 : _T_698; // @[Lookup.scala 33:37]
  assign _T_700 = _T_45 ? 1'h0 : _T_699; // @[Lookup.scala 33:37]
  assign _T_701 = _T_43 ? 1'h0 : _T_700; // @[Lookup.scala 33:37]
  assign _T_702 = _T_41 ? 1'h0 : _T_701; // @[Lookup.scala 33:37]
  assign _T_703 = _T_39 ? 1'h0 : _T_702; // @[Lookup.scala 33:37]
  assign _T_704 = _T_37 ? 1'h0 : _T_703; // @[Lookup.scala 33:37]
  assign _T_705 = _T_35 ? 1'h0 : _T_704; // @[Lookup.scala 33:37]
  assign _T_706 = _T_33 ? 1'h0 : _T_705; // @[Lookup.scala 33:37]
  assign _T_707 = _T_31 ? 1'h0 : _T_706; // @[Lookup.scala 33:37]
  assign _T_708 = _T_29 ? 1'h0 : _T_707; // @[Lookup.scala 33:37]
  assign _T_709 = _T_27 ? 1'h0 : _T_708; // @[Lookup.scala 33:37]
  assign _T_710 = _T_25 ? 1'h0 : _T_709; // @[Lookup.scala 33:37]
  assign _T_711 = _T_23 ? 1'h0 : _T_710; // @[Lookup.scala 33:37]
  assign _T_712 = _T_21 ? 1'h0 : _T_711; // @[Lookup.scala 33:37]
  assign _T_713 = _T_19 ? 1'h0 : _T_712; // @[Lookup.scala 33:37]
  assign _T_714 = _T_17 ? 1'h0 : _T_713; // @[Lookup.scala 33:37]
  assign _T_715 = _T_15 ? 1'h0 : _T_714; // @[Lookup.scala 33:37]
  assign _T_716 = _T_13 ? 1'h0 : _T_715; // @[Lookup.scala 33:37]
  assign _T_717 = _T_11 ? 1'h0 : _T_716; // @[Lookup.scala 33:37]
  assign _T_718 = _T_9 ? 1'h0 : _T_717; // @[Lookup.scala 33:37]
  assign _T_719 = _T_7 ? 1'h0 : _T_718; // @[Lookup.scala 33:37]
  assign _T_720 = _T_5 ? 1'h0 : _T_719; // @[Lookup.scala 33:37]
  assign _T_721 = _T_3 ? 1'h0 : _T_720; // @[Lookup.scala 33:37]
  assign io_pc_sel = _T_1 ? 2'h0 : _T_145; // @[Control.scala 149:16]
  assign io_inst_kill = _T_1 ? 1'h0 : _T_433; // @[Control.scala 150:16]
  assign io_A_sel = _T_1 ? 1'h0 : _T_193; // @[Control.scala 153:14]
  assign io_B_sel = _T_1 ? 1'h0 : _T_241; // @[Control.scala 154:14]
  assign io_imm_sel = _T_1 ? 3'h3 : _T_289; // @[Control.scala 155:14]
  assign io_alu_op = _T_1 ? 4'hb : _T_337; // @[Control.scala 156:14]
  assign io_br_type = _T_1 ? 3'h0 : _T_385; // @[Control.scala 157:14]
  assign io_st_type = _T_1 ? 2'h0 : _T_481; // @[Control.scala 158:14]
  assign io_ld_type = _T_1 ? 3'h0 : _T_529; // @[Control.scala 161:14]
  assign io_wb_sel = _T_1 ? 2'h0 : _T_577; // @[Control.scala 162:14]
  assign io_wb_en = _T_1 | _T_625; // @[Control.scala 163:14]
  assign io_csr_cmd = _T_1 ? 3'h0 : _T_673; // @[Control.scala 164:14]
  assign io_illegal = _T_1 ? 1'h0 : _T_721; // @[Control.scala 165:14]
endmodule
